
module new();
endmodule
