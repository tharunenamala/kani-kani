o "em undi  le"
